
module rf(Clk,WrEn,Ra,Rb,Rw,busW,busA,busB);//que shao R
	input Clk;
	input WrEn;
	input [4:0]Ra,Rb,Rw;
	input [31:0]busW;
	output [31:0]busA,busB;
	
	reg [31:0] R[0:31];

	initial begin
		R[8] = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
		R[9] = 32'b0000_0000_0000_0000_0000_0000_0000_0010;

		R[12] = 32'b0000_0000_0000_0000_0000_0000_0010_0000;
		R[13] = 32'b0000_0000_0000_0000_0000_0000_0010_0000;

		R[15] = 32'b0000_0000_0000_0000_0011_0000_0000_0001;
		R[16] = 32'b0000_0000_0000_0000_0110_0000_0000_0010;

		R[18] = 32'b0000_0000_0000_1010_0000_0000_0000_0001;
		R[19] = 32'b0000_0000_0000_1001_0000_0000_0000_0010;

		R[21] = 32'b0000_0000_0010_0000_0000_0000_0000_0001;
		R[22] = 32'b0000_0000_0100_0000_0000_0000_0000_0010;
	end
	always @(posedge Clk)	begin
		if(WrEn) R[Rw] <= busW;	
		$display(R[10]);
	end

	assign busA = (Ra != 0)? R[Ra]:0;
	assign busB = (Rb != 0)? R[Rb]:0;
endmodule 
